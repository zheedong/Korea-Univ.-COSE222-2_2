/* ********************************************
 *	COSE222 Lab #2
 *
 *	Module: ALU (alu.sv)
 *  - 64-bit 2 input and 1 output ports
 *
 *  Author: Gunjae Koo (gunjaekoo@korea.ac.kr)
 *
 * ********************************************
 */

`timescale 1ns/1ps
`define FF 1    // Flip-flop delay for just better waveform view

module alu
#(  parameter REG_WIDTH = 64 )  // ALU input data width is equal to the width of register file
(
    input   logic [REG_WIDTH-1:0] in1,    // Operand 1
    input   logic [REG_WIDTH-1:0] in2,    // Operand 2
    input   logic [3:0]   alu_control,    // ALU control signal
    output  logic [REG_WIDTH-1:0] result, // ALU output
    output  logic         zero            // Zero detection
);

    always_comb begin
        case (alu_control)
            4'b0010: result = in1 + in2;
            4'b0110: result = in1 - in2;
            4'b0000: result = in1 & in2;
            4'b0001: result = in1 | in2;
            default: result = 0;
		endcase
    end

    assign zero = (result == 0);


endmodule